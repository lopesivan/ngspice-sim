* exemplo 3

v1 1 0 150V
r1 1 2 20
r2 2 0 10
r3 2 3 15
v2 3 0 100V

.op
.END
