How to access parameter values in transient simulation and interactive interpreter

C1 1 0 3uF
R1 1 0 1MEG
V1 1 0 10
.tran 1u 100u

.control
    listing e
    let foo = 123
    define bar(x) ( (x) / foo )
    run
    print foo
    print $&foo  $ print 123
    print bar(12)
    plot V(1)*foo
.endc

.end
