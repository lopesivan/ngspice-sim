How to access parameter values in transient simulation and interactive interpreter

C1 1 0 3uF
R1 1 0 1MEG
V1 1 0 10
.tran 1u 100u

.control
    listing e
    set foo = 123  $ create a new variable
    print $foo     $ prints "123 = 1.230000e+02"
    echo $foo
    define bar(x) ( (x) / $foo )
    tran 1u $foo
    run
    print bar(12)
    plot V(1)*$foo
.endc

.end
