
.TITLE DIODE test

v1 1 0  dc=5
r1 1 2  1k
d1 2 0  D1N750
.model d1n750 D(Vj=.75 Cjo=175p Rs=.25 Eg=1.11 M=.5516 Nbv=1.6989 N=1 Bv=8.1 Fc=.5 Ikf=0 Ibv=20.245m Is=880.5E-18  Xti=3)
.save all @d1[id] @R1[p]

.dc v1 -5 2 0.05

* Control Statements
.control
  run
  plot '-i(v1)' vs v(1)
  plot @d1[id] vs v(1)
  settype power @r1[p]
  plot @r1[p] vs v(1)
.endc

.end
