*SPICE circuit <03468.eps> from XCircuit v3.20
D1 1 5 DI1N4004
V1 5 0 0
D2 1 3 Da1N4004
V2 3 0 0
D3 1 4 Default
V3 4 0 0
V4 1 0 1
.DC V4 0 1400mV 0.2m
.model Da1N4004 D (IS=18.8n RS=0      BV=400 IBV=5.00u CJO=30
+M=0.333   N=2.0  TT=0)
.MODEL DI1N4004 D (IS=76.9n RS=42.0m  BV=400 IBV=5.00u CJO=39.8p
+M=0.333 N=1.45 TT=4.32u)
.MODEL Default D
.end
