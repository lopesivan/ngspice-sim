How to access parameter values in transient simulation and interactive interpreter

.csparam aap = 3
* .param pp = 3*aap
.func omega(x) { 2*aap*x }
* C1 1 0 { aap }
R1 1 0 1MEG
* B1 1 0 I = 25 * aap
* .tran {1u/aap)} {1/aap}
.tran 1u 100u

.control
    listing e
    define bar(x) ( x / aap )
*   tran 1u aap 
    run
    print aap 
    print omega(101)
    run
    plot V(1)*aap
.endc

.end
